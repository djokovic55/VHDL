----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 10/31/2021 09:07:01 AM
-- Design Name: 
-- Module Name: pipo - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity pipo is
    generic(width : positive := 5);
    Port ( 
           d : in STD_LOGIC_VECTOR(width-1 downto 0);
           q : out STD_LOGIC_VECTOR(width-1 downto 0);
           clk : in STD_LOGIC);
end pipo;

architecture Behavioral of pipo is

begin

    process (clk) is 
    begin 
    
        if (rising_edge(clk)) then
            q <= d;
        end if;
        
    end process;
end Behavioral;
